module control_circuit (input clk, input reset, input [5:0] opcode, input [5:0] funct, 
                        output reg IorD, output reg memRead, output reg IRWrite, output reg regDest, output reg regWrite,
                        output reg aluSrcA, output reg [1:0] aluSrcB, output reg [1:0] aluOp, output reg hiWrite,
                        output reg loWrite, output reg [1:0] memToReg, output reg [1:0] pcSrc, output reg pcWrite,output reg branch );

    reg [3:0] state;
    always@(negedge clk)
    begin
        case(state)
        4'b0000 :
        begin
            state=4'b0001;
            IorD=1'b0;
            memRead=1'b1;
            IRWrite=1'b1;
            regDest=1'b0;
            regWrite=1'b0;
            aluSrcA=1'b0;
            aluSrcB=2'b01;
            aluOp=2'b00;
            hiWrite=1'b0;
            loWrite=1'b0;
            memToReg=2'b00;
            pcSrc=2'b10;
            pcWrite=1'b1;
            branch=1'b0;
        end
        4'b0001 :
        begin
            state=4'b0010;
            IorD=1'b0;
            memRead=1'b0;
            IRWrite=1'b0;
            regDest=1'b0;
            regWrite=1'b0;
            aluSrcA=1'b0;
            aluSrcB=2'b11;
            aluOp=2'b00;
            hiWrite=1'b0;
            loWrite=1'b0;
            memToReg=2'b00;
            pcSrc=2'b00;
            pcWrite=1'b0;
            branch=1'b0;
        end
        4'b0010 :
        begin
            case(opcode)
                6'b011000:
                begin
                    state=4'b0100;
                    IorD=1'b0;
                    memRead=1'b0;
                    IRWrite=1'b0;
                    regDest=1'b0;
                    regWrite=1'b0;
                    aluSrcA=1'b1;
                    aluSrcB=2'b00;
                    aluOp=2'b10;
                    hiWrite=1'b0;
                    loWrite=1'b0;
                    memToReg=2'b00;
                    pcSrc=2'b00;
                    pcWrite=1'b0;
                    branch=1'b0;
                end
                6'b010000:
                begin
                    state=4'b0101;
                    IorD=1'b0;
                    memRead=1'b0;
                    IRWrite=1'b0;
                    regDest=1'b1;
                    regWrite=1'b1;
                    aluSrcA=1'b0;
                    aluSrcB=2'b00;
                    aluOp=2'b00;
                    hiWrite=1'b0;
                    loWrite=1'b0;
                    memToReg=2'b01;
                    pcSrc=2'b00;
                    pcWrite=1'b0;
                    branch=1'b0;         
                end
                6'b000100:
                begin
                    state=4'b1000;
                    IorD=1'b0;
                    memRead=1'b0;
                    IRWrite=1'b0;
                    regDest=1'b0;
                    regWrite=1'b0;
                    aluSrcA=1'b1;
                    aluSrcB=2'b00;
                    aluOp=2'b01;
                    hiWrite=1'b0;
                    loWrite=1'b0;
                    memToReg=2'b00;
                    pcSrc=2'b00;
                    pcWrite=1'b0;
                    branch=1'b1;     
                end
                6'b001000:
                begin
                    state=4'b0011;
                        IorD=1'b0;
                        memRead=1'b0;
                        IRWrite=1'b0;
                        regDest=1'b0;
                        regWrite=1'b0;
                        aluSrcA=1'b1;
                        aluSrcB=2'b10;
                        aluOp=2'b00;
                        hiWrite=1'b0;
                        loWrite=1'b0;
                        memToReg=2'b00;
                        pcSrc=2'b00;
                        pcWrite=1'b0;
                        branch=1'b0;     
                end
                6'b100011:
                begin
                    state=4'b0110;
                    IorD=1'b0;
                    memRead=1'b0;
                    IRWrite=1'b0;
                    regDest=1'b0;
                    regWrite=1'b0;
                    aluSrcA=1'b1;
                    aluSrcB=2'b10;
                    aluOp=2'b00;
                    hiWrite=1'b0;
                    loWrite=1'b0;
                    memToReg=2'b00;
                    pcSrc=2'b00;
                    pcWrite=1'b0;
                    branch=1'b0;     
                end
                6'b000010:
                begin
                    state = 4'b0111;
                    IorD=1'b0;
                    memRead=1'b0;
                    IRWrite=1'b0;
                    regDest=1'b0;
                    regWrite=1'b0;
                    aluSrcA=1'b0;
                    aluSrcB=2'b00;
                    aluOp=2'b00;
                    hiWrite=1'b0;
                    loWrite=1'b0;
                    memToReg=2'b00;
                    pcSrc=2'b01;
                    pcWrite=1'b1;
                    branch=1'b0;
                end
                endcase
        end
        4'b0011 :
        begin
            state=4'b1001;
            IorD=1'b0;
            memRead=1'b0;
            IRWrite=1'b0;
            regDest=1'b0;
            regWrite=1'b1;
            aluSrcA=1'b0;
            aluSrcB=2'b00;
            aluOp=2'b00;
            hiWrite=1'b0;
            loWrite=1'b0;
            memToReg=2'b10;
            pcSrc=2'b00;
            pcWrite=1'b0;
            branch=1'b0;
        end
        4'b0100 :
        begin
            state=4'b1010;
            IorD=1'b0;
            memRead=1'b0;
            IRWrite=1'b0;
            regDest=1'b0;
            regWrite=1'b0;
            aluSrcA=1'b0;
            aluSrcB=2'b00;
            aluOp=2'b00;
            hiWrite=1'b1;
            loWrite=1'b1;
            memToReg=2'b00;
            pcSrc=2'b00;
            pcWrite=1'b0;
            branch=1'b0;
        end
        4'b0101 :
        begin
            state=4'b0001;
            IorD=1'b0;
            memRead=1'b1;
            IRWrite=1'b1;
            regDest=1'b0;
            regWrite=1'b0;
            aluSrcA=1'b0;
            aluSrcB=2'b01;
            aluOp=2'b00;
            hiWrite=1'b0;
            loWrite=1'b0;
            memToReg=2'b00;
            pcSrc=2'b10;
            pcWrite=1'b1;
            branch=1'b0;
        end
        4'b0110 :
        begin
            state=4'b1011;
            IorD=1'b1;
                memRead=1'b1;
                IRWrite=1'b0;
                regDest=1'b0;
                regWrite=1'b0;
                aluSrcA=1'b0;
                aluSrcB=2'b00;
                aluOp=2'b00;
                hiWrite=1'b0;
                loWrite=1'b0;
                memToReg=2'b00;
                pcSrc=2'b00;
                pcWrite=1'b0;
                branch=1'b0;
        end
        4'b0111 :
        begin
            state=4'b0001;
            IorD=1'b0;
            memRead=1'b1;
            IRWrite=1'b1;
            regDest=1'b0;
            regWrite=1'b0;
            aluSrcA=1'b0;
            aluSrcB=2'b01;
            aluOp=2'b00;
            hiWrite=1'b0;
            loWrite=1'b0;
            memToReg=2'b00;
            pcSrc=2'b10;
            pcWrite=1'b1;
            branch=1'b0;
        end
        4'b1000 :
        begin
            state=4'b0001;
            IorD=1'b0;
            memRead=1'b1;
            IRWrite=1'b1;
            regDest=1'b0;
            regWrite=1'b0;
            aluSrcA=1'b0;
            aluSrcB=2'b01;
            aluOp=2'b00;
            hiWrite=1'b0;
            loWrite=1'b0;
            memToReg=2'b00;
            pcSrc=2'b10;
            pcWrite=1'b1;
            branch=1'b0;
        end
        4'b1001 :
        begin
            state=4'b0001;
            IorD=1'b0;
            memRead=1'b1;
            IRWrite=1'b1;
            regDest=1'b0;
            regWrite=1'b0;
            aluSrcA=1'b0;
            aluSrcB=2'b01;
            aluOp=2'b00;
            hiWrite=1'b0;
            loWrite=1'b0;
            memToReg=2'b00;
            pcSrc=2'b10;
            pcWrite=1'b1;
            branch=1'b0;
        end
        4'b1010 :
        begin
            state=4'b0001;
            IorD=1'b0;
            memRead=1'b1;
            IRWrite=1'b1;
            regDest=1'b0;
            regWrite=1'b0;
            aluSrcA=1'b0;
            aluSrcB=2'b01;
            aluOp=2'b00;
            hiWrite=1'b0;
            loWrite=1'b0;
            memToReg=2'b00;
            pcSrc=2'b10;
            pcWrite=1'b1;
            branch=1'b0; 
        end
        4'b1011 :
        begin
                state=4'b1100;
                IorD=1'b0;
                memRead=1'b0;
                IRWrite=1'b0;
                regDest=1'b0;
                regWrite=1'b1;
                aluSrcA=1'b0;
                aluSrcB=2'b00;
                aluOp=2'b00;
                hiWrite=1'b0;
                loWrite=1'b0;
                memToReg=2'b00;
                pcSrc=2'b00;
                pcWrite=1'b0;
                branch=1'b0;
        end
        4'b1100 :
        begin
            state=4'b0001;
            IorD=1'b0;
            memRead=1'b1;
            IRWrite=1'b1;
            regDest=1'b0;
            regWrite=1'b0;
            aluSrcA=1'b0;
            aluSrcB=2'b01;
            aluOp=2'b00;
            hiWrite=1'b0;
            loWrite=1'b0;
            memToReg=2'b00;
            pcSrc=2'b10;
            pcWrite=1'b1;
            branch=1'b0;
        end
        default:
        begin
            state=4'b0000;
            IorD=1'b0;
            memRead=1'b0;
            IRWrite=1'b0;
            regDest=1'b0;
            regWrite=1'b0;
            aluSrcA=1'b0;
            aluSrcB=2'b00;
            aluOp=2'b00;
            hiWrite=1'b0;
            loWrite=1'b0;
            memToReg=2'b00;
            pcSrc=2'b11;
            pcWrite=1'b0;
            branch=1'b0;
        end
        endcase
    end



endmodule